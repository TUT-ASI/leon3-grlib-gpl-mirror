-- High Speed Serial Links
  constant CFG_HSSL_EN   : integer := CONFIG_GRHSSL_ENABLE;
  constant CFG_HSSL_NUM  : integer := CONFIG_GRHSSL_NUM;
  constant CFG_HSSL_SPFI : integer := CONFIG_GRHSSL_SPFI;
  constant CFG_HSSL_WIZL : integer := CONFIG_GRHSSL_WIZL;
