
package version is
  constant grlib_version : integer := 2020200;
  constant grlib_build : integer := 4254;
end;
