-- GRDMAC2 interface
  constant CFG_GRDMAC2       : integer := CONFIG_GRDMAC2_ENABLE;
  constant CFG_GRDMAC2ACC    : integer := CONFIG_GRDMAC2ACC;
  constant CFG_GRDMAC2FT     : integer := CONFIG_GRDMAC2FT;
  constant CFG_GRDMAC2ABITS  : integer := CONFIG_GRDMAC2ABITS;
  constant CFG_GRDMAC2DBITS  : integer := CONFIG_GRDMAC2DBITS;
  
