-- SPI controller
  constant CFG_SPICTRL_ENABLE : integer := CONFIG_SPICTRL_ENABLE;
  constant CFG_SPICTRL_SLVS   : integer := CONFIG_SPICTRL_SLVS;
  constant CFG_SPICTRL_FIFO   : integer := CONFIG_SPICTRL_FIFO;
  constant CFG_SPICTRL_SLVREG : integer := CONFIG_SPICTRL_SLVREG;
  constant CFG_SPICTRL_ODMODE : integer := CONFIG_SPICTRL_ODMODE;
  constant CFG_SPICTRL_AM     : integer := CONFIG_SPICTRL_AM;
  constant CFG_SPICTRL_ASEL   : integer := CONFIG_SPICTRL_ASEL;

