package rev is
  constant REVISION : integer := 130;
end;
