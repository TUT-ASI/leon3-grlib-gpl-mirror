package rev is
  constant REVISION : integer := 140;
end;
