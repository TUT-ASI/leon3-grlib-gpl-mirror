
package version is
  constant grlib_version : integer := 2020400;
  constant grlib_build : integer := 4261;
end;
