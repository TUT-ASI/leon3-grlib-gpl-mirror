package rev is
  constant REVISION : integer := 120;
end;
