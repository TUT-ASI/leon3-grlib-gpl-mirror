--LEON5 processor system
  constant CFG_NCPU    : integer := CONFIG_PROC_NUM;
  constant CFG_FPUTYPE : integer := CONFIG_FPU;
  constant CFG_AHBW    : integer := CONFIG_AHBW;
  constant CFG_BWMASK  : integer := 16#CONFIG_BWMASK#;
  constant CFG_DFIXED  : integer := 16#CONFIG_CACHE_FIXED#;

