-- LEON3 Statistics Module
  constant CFG_L3S_ENABLE   : integer := CONFIG_L3S_ENABLE;
  constant CFG_L3S_CNT      : integer := CONFIG_L3S_CNT;
  constant CFG_L3S_NMAX     : integer := CONFIG_L3S_NMAX;

