
package version is
  constant grlib_version : integer := 2024200;
  constant grlib_build : integer := 4293;
end;
