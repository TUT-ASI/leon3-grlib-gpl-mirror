-- HPS
  constant CFG_HPS2FPGA   : integer := CONFIG_HPS2FPGA;
  constant CFG_FPGA2HPS   : integer := CONFIG_FPGA2HPS;
  constant CFG_HPS_RESET  : integer := CONFIG_HPS_RESET;

