-- USB Host Controller
  constant CFG_USBHC          : integer := CONFIG_GRUSBHC_ENABLE;
  constant CFG_USBHC_NPORTS   : integer := CONFIG_GRUSBHC_NPORTS;
  constant CFG_USBHC_EHC      : integer := CONFIG_GRUSBHC_EHC;
  constant CFG_USBHC_UHC      : integer := CONFIG_GRUSBHC_UHC;
  constant CFG_USBHC_NCC      : integer := CONFIG_GRUSBHC_NCC;
  constant CFG_USBHC_NPCC     : integer := CONFIG_GRUSBHC_NPCC;
  constant CFG_USBHC_PRR      : integer := CONFIG_GRUSBHC_PRR;
  constant CFG_USBHC_PR1      : integer := CONFIG_GRUSBHC_PORTROUTE1;
  constant CFG_USBHC_PR2      : integer := CONFIG_GRUSBHC_PORTROUTE2;
  constant CFG_USBHC_ENDIAN   : integer := CONFIG_GRUSBHC_ENDIAN;
  constant CFG_USBHC_BEREGS   : integer := CONFIG_GRUSBHC_BEREGS;
  constant CFG_USBHC_BEDESC   : integer := CONFIG_GRUSBHC_BEDESC;
  constant CFG_USBHC_BLO      : integer := CONFIG_GRUSBHC_BLO;
  constant CFG_USBHC_BWRD     : integer := CONFIG_GRUSBHC_BWRD;
  constant CFG_USBHC_UTM      : integer := CONFIG_GRUSBHC_UTMTYPE;
  constant CFG_USBHC_VBUSCONF : integer := CONFIG_GRUSBHC_VBUSCONF;

