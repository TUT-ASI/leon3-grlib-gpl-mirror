package rev is
  constant REVISION : integer := 100;
end;
