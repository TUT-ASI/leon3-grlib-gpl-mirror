-- megafunction wizard: %Triple-Speed Ethernet v13.1%
-- GENERATION: XML
-- sgmii2gmii.vhd

-- Generated using ACDS version 13.1 162 at 2013.11.29.14:56:05

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sgmii2gmii is
	port (
		ref_clk        : in  std_logic                     := '0';             --  pcs_ref_clk_clock_connection.clk
		clk            : in  std_logic                     := '0';             -- control_port_clock_connection.clk
		reset          : in  std_logic                     := '0';             --              reset_connection.reset
		address        : in  std_logic_vector(4 downto 0)  := (others => '0'); --                  control_port.address
		readdata       : out std_logic_vector(15 downto 0);                    --                              .readdata
		read           : in  std_logic                     := '0';             --                              .read
		writedata      : in  std_logic_vector(15 downto 0) := (others => '0'); --                              .writedata
		write          : in  std_logic                     := '0';             --                              .write
		waitrequest    : out std_logic;                                        --                              .waitrequest
		tx_clk         : out std_logic;                                        -- pcs_transmit_clock_connection.clk
		rx_clk         : out std_logic;                                        --  pcs_receive_clock_connection.clk
		reset_tx_clk   : in  std_logic                     := '0';             -- pcs_transmit_reset_connection.reset
		reset_rx_clk   : in  std_logic                     := '0';             --  pcs_receive_reset_connection.reset
		gmii_rx_dv     : out std_logic;                                        --               gmii_connection.gmii_rx_dv
		gmii_rx_d      : out std_logic_vector(7 downto 0);                     --                              .gmii_rx_d
		gmii_rx_err    : out std_logic;                                        --                              .gmii_rx_err
		gmii_tx_en     : in  std_logic                     := '0';             --                              .gmii_tx_en
		gmii_tx_d      : in  std_logic_vector(7 downto 0)  := (others => '0'); --                              .gmii_tx_d
		gmii_tx_err    : in  std_logic                     := '0';             --                              .gmii_tx_err
		tx_clkena      : out std_logic;                                        --       clock_enable_connection.tx_clkena
		rx_clkena      : out std_logic;                                        --                              .rx_clkena
		mii_rx_dv      : out std_logic;                                        --                mii_connection.mii_rx_dv
		mii_rx_d       : out std_logic_vector(3 downto 0);                     --                              .mii_rx_d
		mii_rx_err     : out std_logic;                                        --                              .mii_rx_err
		mii_tx_en      : in  std_logic                     := '0';             --                              .mii_tx_en
		mii_tx_d       : in  std_logic_vector(3 downto 0)  := (others => '0'); --                              .mii_tx_d
		mii_tx_err     : in  std_logic                     := '0';             --                              .mii_tx_err
		mii_col        : out std_logic;                                        --                              .mii_col
		mii_crs        : out std_logic;                                        --                              .mii_crs
		set_10         : out std_logic;                                        --       sgmii_status_connection.set_10
		set_1000       : out std_logic;                                        --                              .set_1000
		set_100        : out std_logic;                                        --                              .set_100
		hd_ena         : out std_logic;                                        --                              .hd_ena
		led_crs        : out std_logic;                                        --         status_led_connection.crs
		led_link       : out std_logic;                                        --                              .link
		led_col        : out std_logic;                                        --                              .col
		led_an         : out std_logic;                                        --                              .an
		led_char_err   : out std_logic;                                        --                              .char_err
		led_disp_err   : out std_logic;                                        --                              .disp_err
		rx_recovclkout : out std_logic;                                        --     serdes_control_connection.export
		txp            : out std_logic;                                        --             serial_connection.txp
		rxp            : in  std_logic                     := '0'              --                              .rxp
	);
end entity sgmii2gmii;

architecture rtl of sgmii2gmii is
	component sgmii2gmii_0002 is
		port (
			ref_clk        : in  std_logic                     := 'X';             -- clk
			clk            : in  std_logic                     := 'X';             -- clk
			reset          : in  std_logic                     := 'X';             -- reset
			address        : in  std_logic_vector(4 downto 0)  := (others => 'X'); -- address
			readdata       : out std_logic_vector(15 downto 0);                    -- readdata
			read           : in  std_logic                     := 'X';             -- read
			writedata      : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			write          : in  std_logic                     := 'X';             -- write
			waitrequest    : out std_logic;                                        -- waitrequest
			tx_clk         : out std_logic;                                        -- clk
			rx_clk         : out std_logic;                                        -- clk
			reset_tx_clk   : in  std_logic                     := 'X';             -- reset
			reset_rx_clk   : in  std_logic                     := 'X';             -- reset
			gmii_rx_dv     : out std_logic;                                        -- gmii_rx_dv
			gmii_rx_d      : out std_logic_vector(7 downto 0);                     -- gmii_rx_d
			gmii_rx_err    : out std_logic;                                        -- gmii_rx_err
			gmii_tx_en     : in  std_logic                     := 'X';             -- gmii_tx_en
			gmii_tx_d      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- gmii_tx_d
			gmii_tx_err    : in  std_logic                     := 'X';             -- gmii_tx_err
			tx_clkena      : out std_logic;                                        -- tx_clkena
			rx_clkena      : out std_logic;                                        -- rx_clkena
			mii_rx_dv      : out std_logic;                                        -- mii_rx_dv
			mii_rx_d       : out std_logic_vector(3 downto 0);                     -- mii_rx_d
			mii_rx_err     : out std_logic;                                        -- mii_rx_err
			mii_tx_en      : in  std_logic                     := 'X';             -- mii_tx_en
			mii_tx_d       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- mii_tx_d
			mii_tx_err     : in  std_logic                     := 'X';             -- mii_tx_err
			mii_col        : out std_logic;                                        -- mii_col
			mii_crs        : out std_logic;                                        -- mii_crs
			set_10         : out std_logic;                                        -- set_10
			set_1000       : out std_logic;                                        -- set_1000
			set_100        : out std_logic;                                        -- set_100
			hd_ena         : out std_logic;                                        -- hd_ena
			led_crs        : out std_logic;                                        -- crs
			led_link       : out std_logic;                                        -- link
			led_col        : out std_logic;                                        -- col
			led_an         : out std_logic;                                        -- an
			led_char_err   : out std_logic;                                        -- char_err
			led_disp_err   : out std_logic;                                        -- disp_err
			rx_recovclkout : out std_logic;                                        -- export
			txp            : out std_logic;                                        -- txp
			rxp            : in  std_logic                     := 'X'              -- rxp
		);
	end component sgmii2gmii_0002;

begin

	sgmii2gmii_inst : component sgmii2gmii_0002
		port map (
			ref_clk        => ref_clk,        --  pcs_ref_clk_clock_connection.clk
			clk            => clk,            -- control_port_clock_connection.clk
			reset          => reset,          --              reset_connection.reset
			address        => address,        --                  control_port.address
			readdata       => readdata,       --                              .readdata
			read           => read,           --                              .read
			writedata      => writedata,      --                              .writedata
			write          => write,          --                              .write
			waitrequest    => waitrequest,    --                              .waitrequest
			tx_clk         => tx_clk,         -- pcs_transmit_clock_connection.clk
			rx_clk         => rx_clk,         --  pcs_receive_clock_connection.clk
			reset_tx_clk   => reset_tx_clk,   -- pcs_transmit_reset_connection.reset
			reset_rx_clk   => reset_rx_clk,   --  pcs_receive_reset_connection.reset
			gmii_rx_dv     => gmii_rx_dv,     --               gmii_connection.gmii_rx_dv
			gmii_rx_d      => gmii_rx_d,      --                              .gmii_rx_d
			gmii_rx_err    => gmii_rx_err,    --                              .gmii_rx_err
			gmii_tx_en     => gmii_tx_en,     --                              .gmii_tx_en
			gmii_tx_d      => gmii_tx_d,      --                              .gmii_tx_d
			gmii_tx_err    => gmii_tx_err,    --                              .gmii_tx_err
			tx_clkena      => tx_clkena,      --       clock_enable_connection.tx_clkena
			rx_clkena      => rx_clkena,      --                              .rx_clkena
			mii_rx_dv      => mii_rx_dv,      --                mii_connection.mii_rx_dv
			mii_rx_d       => mii_rx_d,       --                              .mii_rx_d
			mii_rx_err     => mii_rx_err,     --                              .mii_rx_err
			mii_tx_en      => mii_tx_en,      --                              .mii_tx_en
			mii_tx_d       => mii_tx_d,       --                              .mii_tx_d
			mii_tx_err     => mii_tx_err,     --                              .mii_tx_err
			mii_col        => mii_col,        --                              .mii_col
			mii_crs        => mii_crs,        --                              .mii_crs
			set_10         => set_10,         --       sgmii_status_connection.set_10
			set_1000       => set_1000,       --                              .set_1000
			set_100        => set_100,        --                              .set_100
			hd_ena         => hd_ena,         --                              .hd_ena
			led_crs        => led_crs,        --         status_led_connection.crs
			led_link       => led_link,       --                              .link
			led_col        => led_col,        --                              .col
			led_an         => led_an,         --                              .an
			led_char_err   => led_char_err,   --                              .char_err
			led_disp_err   => led_disp_err,   --                              .disp_err
			rx_recovclkout => rx_recovclkout, --     serdes_control_connection.export
			txp            => txp,            --             serial_connection.txp
			rxp            => rxp             --                              .rxp
		);

end architecture rtl; -- of sgmii2gmii
-- Retrieval info: <?xml version="1.0"?>
--<!--
--	Generated by Altera MegaWizard Launcher Utility version 1.0
--	************************************************************
--	THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--	************************************************************
--	Copyright (C) 1991-2013 Altera Corporation
--	Any megafunction design, and related net list (encrypted or decrypted),
--	support information, device programming or simulation file, and any other
--	associated documentation or information provided by Altera or a partner
--	under Altera's Megafunction Partnership Program may be used only to
--	program PLD devices (but not masked PLD devices) from Altera.  Any other
--	use of such megafunction design, net list, support information, device
--	programming or simulation file, or any other related documentation or
--	information is prohibited for any other purpose, including, but not
--	limited to modification, reverse engineering, de-compiling, or use with
--	any other silicon devices, unless such use is explicitly licensed under
--	a separate agreement with Altera or a megafunction partner.  Title to
--	the intellectual property, including patents, copyrights, trademarks,
--	trade secrets, or maskworks, embodied in any such megafunction design,
--	net list, support information, device programming or simulation file, or
--	any other related documentation or information provided by Altera or a
--	megafunction partner, remains with Altera, the megafunction partner, or
--	their respective licensors.  No other licenses, including any licenses
--	needed under any third party's intellectual property, are provided herein.
---->
-- Retrieval info: <instance entity-name="altera_eth_tse" version="13.1" >
-- Retrieval info: 	<generic name="deviceFamilyName" value="Stratix IV" />
-- Retrieval info: 	<generic name="core_variation" value="PCS_ONLY" />
-- Retrieval info: 	<generic name="ifGMII" value="MII_GMII" />
-- Retrieval info: 	<generic name="enable_use_internal_fifo" value="true" />
-- Retrieval info: 	<generic name="max_channels" value="1" />
-- Retrieval info: 	<generic name="use_misc_ports" value="true" />
-- Retrieval info: 	<generic name="transceiver_type" value="LVDS_IO" />
-- Retrieval info: 	<generic name="enable_hd_logic" value="true" />
-- Retrieval info: 	<generic name="enable_gmii_loopback" value="false" />
-- Retrieval info: 	<generic name="enable_sup_addr" value="false" />
-- Retrieval info: 	<generic name="stat_cnt_ena" value="true" />
-- Retrieval info: 	<generic name="ext_stat_cnt_ena" value="false" />
-- Retrieval info: 	<generic name="ena_hash" value="false" />
-- Retrieval info: 	<generic name="enable_shift16" value="true" />
-- Retrieval info: 	<generic name="enable_mac_flow_ctrl" value="false" />
-- Retrieval info: 	<generic name="enable_mac_vlan" value="false" />
-- Retrieval info: 	<generic name="enable_magic_detect" value="true" />
-- Retrieval info: 	<generic name="useMDIO" value="false" />
-- Retrieval info: 	<generic name="mdio_clk_div" value="40" />
-- Retrieval info: 	<generic name="enable_ena" value="32" />
-- Retrieval info: 	<generic name="eg_addr" value="11" />
-- Retrieval info: 	<generic name="ing_addr" value="11" />
-- Retrieval info: 	<generic name="phy_identifier" value="0" />
-- Retrieval info: 	<generic name="enable_sgmii" value="true" />
-- Retrieval info: 	<generic name="export_pwrdn" value="false" />
-- Retrieval info: 	<generic name="enable_alt_reconfig" value="false" />
-- Retrieval info: 	<generic name="starting_channel_number" value="0" />
-- Retrieval info: 	<generic name="phyip_pll_type" value="CMU" />
-- Retrieval info: 	<generic name="phyip_en_synce_support" value="false" />
-- Retrieval info: 	<generic name="phyip_pma_bonding_mode" value="x1" />
-- Retrieval info: 	<generic name="nf_phyip_rcfg_enable" value="false" />
-- Retrieval info: 	<generic name="enable_timestamping" value="false" />
-- Retrieval info: 	<generic name="enable_ptp_1step" value="false" />
-- Retrieval info: 	<generic name="tstamp_fp_width" value="4" />
-- Retrieval info: 	<generic name="AUTO_DEVICE" value="Unknown" />
-- Retrieval info: </instance>
-- IPFS_FILES : sgmii2gmii.vho
-- RELATED_FILES: sgmii2gmii.vhd, sgmii2gmii_0002.v, altera_eth_tse_pcs_pma_lvds.v, altera_tse_align_sync.v, altera_tse_dec10b8b.v, altera_tse_dec_func.v, altera_tse_enc8b10b.v, altera_tse_top_autoneg.v, altera_tse_carrier_sense.v, altera_tse_clk_gen.v, altera_tse_sgmii_clk_div.v, altera_tse_sgmii_clk_enable.v, altera_tse_rx_encapsulation.v, altera_tse_tx_encapsulation.v, altera_tse_rx_encapsulation_strx_gx.v, altera_tse_pcs_control.v, altera_tse_pcs_host_control.v, altera_tse_mdio_reg.v, altera_tse_mii_rx_if_pcs.v, altera_tse_mii_tx_if_pcs.v, altera_tse_rx_sync.v, altera_tse_sgmii_clk_cntl.v, altera_tse_colision_detect.v, altera_tse_rx_converter.v, altera_tse_rx_fifo_rd.v, altera_tse_top_rx_converter.v, altera_tse_top_sgmii.v, altera_tse_top_sgmii_strx_gx.v, altera_tse_top_tx_converter.v, altera_tse_tx_converter.v, altera_tse_top_1000_base_x.v, altera_tse_top_1000_base_x_strx_gx.v, altera_tse_top_pcs.v, altera_tse_top_pcs_strx_gx.v, altera_tse_top_rx.v, altera_tse_top_tx.v, altera_tse_lvds_reset_sequencer.v, altera_tse_lvds_reverse_loopback.v, altera_tse_pma_lvds_rx_av.v, altera_tse_pma_lvds_rx.v, altera_tse_pma_lvds_tx.v, altera_tse_false_path_marker.v, altera_tse_reset_synchronizer.v, altera_tse_clock_crosser.v, altera_tse_a_fifo_13.v, altera_tse_a_fifo_24.v, altera_tse_a_fifo_34.v, altera_tse_a_fifo_opt_1246.v, altera_tse_a_fifo_opt_14_44.v, altera_tse_a_fifo_opt_36_10.v, altera_tse_gray_cnt.v, altera_tse_sdpm_altsyncram.v, altera_tse_altsyncram_dpm_fifo.v, altera_tse_bin_cnt.v, altera_tse_ph_calculator.sv, altera_tse_sdpm_gen.v, altera_tse_dc_fifo.v
