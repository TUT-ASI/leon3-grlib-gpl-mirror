
package version is
  constant grlib_version : integer := 2025100;
  constant grlib_build : integer := 4296;
end;
