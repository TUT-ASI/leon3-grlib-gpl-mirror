
package version is
  constant grlib_version : integer := 2022100;
  constant grlib_build : integer := 4272;
end;
