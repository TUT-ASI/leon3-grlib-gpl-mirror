
package version is
  constant grlib_version : integer := 2023100;
  constant grlib_build : integer := 4282;
end;
