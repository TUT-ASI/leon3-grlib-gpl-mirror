
package version is
  constant grlib_version : integer := 2025200;
  constant grlib_build : integer := 4298;
end;
