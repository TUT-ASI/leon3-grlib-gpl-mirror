-- NOEL-V processor core
  constant CFG_NOELV  	        : integer := CONFIG_NOELV;
  constant CFG_NCPU             : integer := CONFIG_PROC_NUM;
  constant CFG_CFG              : integer := CONFIG_PROC_CFG;
  constant CFG_NODBUS           : integer := CONFIG_PROC_NODBUS;
  constant CFG_DISAS            : integer := 3*CONFIG_IU_DISAS;

