
package version is
  constant grlib_version : integer := 2019200;
  constant grlib_build : integer := 4241;
end;
