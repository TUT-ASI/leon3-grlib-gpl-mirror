-- CoreMP7 with GRLIB bridge
  constant CFG_CMP7GRLIB          : integer := CONFIG_CMP7GRLIB;
  constant CFG_CMP7GRLIB_DEBUG    : integer := CONFIG_CMP7GRLIB_DEBUG;
  constant CFG_CMP7GRLIB_SYNCFIQ  : integer := CONFIG_CMP7GRLIB_SYNCFIQ;
  constant CFG_CMP7GRLIB_SYNCIRQ  : integer := CONFIG_CMP7GRLIB_SYNCIRQ;
  
