
package version is
  constant grlib_version : integer := 2018100;
  constant grlib_build : integer := 4217;
end;
