
package version is
  constant grlib_version : integer := 2021200;
  constant grlib_build : integer := 4267;
end;
