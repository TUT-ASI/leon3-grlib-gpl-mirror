package rev is
  constant REVISION : integer := 110;
end;
