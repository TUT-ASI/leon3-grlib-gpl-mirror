
package version is
  constant grlib_version : integer := 2022400;
  constant grlib_build : integer := 4280;
end;
