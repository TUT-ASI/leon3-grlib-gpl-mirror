-- GRCANFD interface
  constant CFG_GRCANFD       : integer := CONFIG_GRCANFD_ENABLE;
  constant CFG_GRCANFDIRQ    : integer := CONFIG_GRCANFDIRQ;
  constant CFG_GRCANFDSINGLE : integer := CONFIG_GRCANFDSINGLE;

