package rev is
  constant REVISION : integer := 111;
end;
