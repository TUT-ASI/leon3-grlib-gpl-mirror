-- pragma translate_off
use std.textio.all;
-- pragma translate_on
package version is
  constant grlib_version : integer := 1307;
-- pragma translate_off
  constant grlib_date : string := "20140416";
-- pragma translate_on
  constant grlib_build : integer := 4144;
end;
