-- pragma translate_off
use std.textio.all;
-- pragma translate_on
package version is
  constant grlib_version : integer := 1300;
-- pragma translate_off
  constant grlib_date : string := "20130724";
-- pragma translate_on
  constant grlib_build : integer := 4133;
end;
