
package version is
  constant grlib_version : integer := 2024400;
  constant grlib_build : integer := 4295;
end;
