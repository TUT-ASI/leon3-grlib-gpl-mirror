-- Version and Revision Register
  constant CFG_GRVERSION_ENABLE : integer := CONFIG_GRVERSION_ENABLE;
  constant CFG_GRVERSION_VERSION  : integer := 16#CONFIG_GRVERSION_VERSION#;
  constant CFG_GRVERSION_REVISION  : integer := 16#CONFIG_GRVERSION_REVISION#;

