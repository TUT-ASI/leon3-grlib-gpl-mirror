
package version is
  constant grlib_version : integer := 2020100;
  constant grlib_build : integer := 4251;
end;
