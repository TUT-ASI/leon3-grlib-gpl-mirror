
package version is
  constant grlib_version : integer := 2022200;
  constant grlib_build : integer := 4274;
end;
