-- Version: 
-- VHDL Black Box file 
-- 

library ieee;
use ieee.std_logic_1164.all;
library smartfusion2;
use smartfusion2.all;

entity SERDESIF_0 is
	generic (
		INIT:std_logic_vector := x"0";
		ACT_CONFIG:string := "";
		ACT_SIM:integer := 0	);
   port( 
       APB_PRDATA : out std_logic_vector(31 downto 0);
       APB_PREADY : out std_logic;
       APB_PSLVERR : out std_logic;
       ATXCLKSTABLE : out std_logic_vector(1 downto 0);
       EPCS_READY : out std_logic_vector(1 downto 0);
       EPCS_RXCLK : out std_logic_vector(1 downto 0);
       EPCS_RXCLK_0 : out std_logic;
       EPCS_RXCLK_1 : out std_logic;
       EPCS_RXDATA : out std_logic_vector(39 downto 0);
       EPCS_RXIDLE : out std_logic_vector(1 downto 0);
       EPCS_RXRSTN : out std_logic_vector(1 downto 0);
       EPCS_RXVAL : out std_logic_vector(1 downto 0);
       EPCS_TXCLK : out std_logic_vector(1 downto 0);
       EPCS_TXCLK_0 : out std_logic;
       EPCS_TXCLK_1 : out std_logic;
       EPCS_TXRSTN : out std_logic_vector(1 downto 0);
       FATC_RESET_N : out std_logic;
       H2FCALIB0 : out std_logic;
       H2FCALIB1 : out std_logic;
       M_ARADDR : out std_logic_vector(31 downto 0);
       M_ARBURST : out std_logic_vector(1 downto 0);
       M_ARID : out std_logic_vector(3 downto 0);
       M_ARLEN : out std_logic_vector(3 downto 0);
       M_ARSIZE : out std_logic_vector(1 downto 0);
       M_ARVALID : out std_logic;
       M_AWADDR_HADDR : out std_logic_vector(31 downto 0);
       M_AWBURST_HTRANS : out std_logic_vector(1 downto 0);
       M_AWID : out std_logic_vector(3 downto 0);
       M_AWLEN_HBURST : out std_logic_vector(3 downto 0);
       M_AWSIZE_HSIZE : out std_logic_vector(1 downto 0);
       M_AWVALID_HWRITE : out std_logic;
       M_BREADY : out std_logic;
       M_RREADY : out std_logic;
       M_WDATA_HWDATA : out std_logic_vector(63 downto 0);
       M_WID : out std_logic_vector(3 downto 0);
       M_WLAST : out std_logic;
       M_WSTRB : out std_logic_vector(7 downto 0);
       M_WVALID : out std_logic;
       PCIE_SYSTEM_INT : out std_logic;
       PLL_LOCK_INT : out std_logic;
       PLL_LOCKLOST_INT : out std_logic;
       S_ARREADY : out std_logic;
       S_AWREADY : out std_logic;
       S_BID : out std_logic_vector(3 downto 0);
       S_BRESP_HRESP : out std_logic_vector(1 downto 0);
       S_BVALID : out std_logic;
       S_RDATA_HRDATA : out std_logic_vector(63 downto 0);
       S_RID : out std_logic_vector(3 downto 0);
       S_RLAST : out std_logic;
       S_RRESP : out std_logic_vector(1 downto 0);
       S_RVALID : out std_logic;
       S_WREADY_HREADYOUT : out std_logic;
       SPLL_LOCK : out std_logic;
       WAKE_N : out std_logic;
       XAUI_OUT_CLK : out std_logic;
       APB_CLK : in std_logic;
       APB_PADDR : in std_logic_vector(13 downto 2);
       APB_PENABLE : in std_logic;
       APB_PSEL : in std_logic;
       APB_PWDATA : in std_logic_vector(31 downto 0);
       APB_PWRITE : in std_logic;
       APB_RSTN : in std_logic;
       CLK_BASE : in std_logic;
       EPCS_PWRDN : in std_logic_vector(1 downto 0);
       EPCS_RSTN : in std_logic_vector(1 downto 0);
       EPCS_RXERR : in std_logic_vector(1 downto 0);
       EPCS_TXDATA : in std_logic_vector(39 downto 0);
       EPCS_TXOOB : in std_logic_vector(1 downto 0);
       EPCS_TXVAL : in std_logic_vector(1 downto 0);
       F2HCALIB0 : in std_logic;
       F2HCALIB1 : in std_logic;
       FAB_PLL_LOCK : in std_logic;
       FAB_REF_CLK : in std_logic;
       M_ARREADY : in std_logic;
       M_AWREADY : in std_logic;
       M_BID : in std_logic_vector(3 downto 0);
       M_BRESP_HRESP : in std_logic_vector(1 downto 0);
       M_BVALID : in std_logic;
       M_RDATA_HRDATA : in std_logic_vector(63 downto 0);
       M_RID : in std_logic_vector(3 downto 0);
       M_RLAST : in std_logic;
       M_RRESP : in std_logic_vector(1 downto 0);
       M_RVALID : in std_logic;
       M_WREADY_HREADY : in std_logic;
       PCIE_INTERRUPT : in std_logic_vector(3 downto 0);
       PERST_N : in std_logic;
       S_ARADDR : in std_logic_vector(31 downto 0);
       S_ARBURST : in std_logic_vector(1 downto 0);
       S_ARID : in std_logic_vector(3 downto 0);
       S_ARLEN : in std_logic_vector(3 downto 0);
       S_ARLOCK : in std_logic_vector(1 downto 0);
       S_ARSIZE : in std_logic_vector(1 downto 0);
       S_ARVALID : in std_logic;
       S_AWADDR_HADDR : in std_logic_vector(31 downto 0);
       S_AWBURST_HTRANS : in std_logic_vector(1 downto 0);
       S_AWID_HSEL : in std_logic_vector(3 downto 0);
       S_AWLEN_HBURST : in std_logic_vector(3 downto 0);
       S_AWLOCK : in std_logic_vector(1 downto 0);
       S_AWSIZE_HSIZE : in std_logic_vector(1 downto 0);
       S_AWVALID_HWRITE : in std_logic;
       S_BREADY_HREADY : in std_logic;
       S_RREADY : in std_logic;
       S_WDATA_HWDATA : in std_logic_vector(63 downto 0);
       S_WID : in std_logic_vector(3 downto 0);
       S_WLAST : in std_logic;
       S_WSTRB : in std_logic_vector(7 downto 0);
       S_WVALID : in std_logic;
       SERDESIF_CORE_RESET_N : in std_logic;
       SERDESIF_PHY_RESET_N : in std_logic;
       WAKE_REQ : in std_logic;
       XAUI_FB_CLK : in std_logic;
       RXD3_P : in std_logic;
       RXD2_P : in std_logic;
       RXD1_P : in std_logic;
       RXD0_P : in std_logic;
       RXD3_N : in std_logic;
       RXD2_N : in std_logic;
       RXD1_N : in std_logic;
       RXD0_N : in std_logic;
       TXD3_P : out std_logic;
       TXD2_P : out std_logic;
       TXD1_P : out std_logic;
       TXD0_P : out std_logic;
       TXD3_N : out std_logic;
       TXD2_N : out std_logic;
       TXD1_N : out std_logic;
       TXD0_N : out std_logic;
       REFCLK0 : in std_logic;
       REFCLK1 : in std_logic
   );
end SERDESIF_0;
architecture DEF_ARCH of SERDESIF_0 is 

   attribute black_box : boolean;
   attribute black_box of DEF_ARCH : architecture is true;
   attribute ment_tsu0: string;
   attribute ment_tsu0 of DEF_ARCH : architecture is " APB_PADDR[10]->APB_CLK=0.085";
   attribute ment_tsu1: string;
   attribute ment_tsu1 of DEF_ARCH : architecture is " APB_PADDR[11]->APB_CLK=-0.125";
   attribute ment_tsu2: string;
   attribute ment_tsu2 of DEF_ARCH : architecture is " APB_PADDR[12]->APB_CLK=1.385";
   attribute ment_tsu3: string;
   attribute ment_tsu3 of DEF_ARCH : architecture is " APB_PADDR[13]->APB_CLK=1.405";
   attribute ment_tsu4: string;
   attribute ment_tsu4 of DEF_ARCH : architecture is " APB_PADDR[2]->APB_CLK=4.043";
   attribute ment_tsu5: string;
   attribute ment_tsu5 of DEF_ARCH : architecture is " APB_PADDR[3]->APB_CLK=4.683";
   attribute ment_tsu6: string;
   attribute ment_tsu6 of DEF_ARCH : architecture is " APB_PADDR[4]->APB_CLK=5.548";
   attribute ment_tsu7: string;
   attribute ment_tsu7 of DEF_ARCH : architecture is " APB_PADDR[5]->APB_CLK=3.703";
   attribute ment_tsu8: string;
   attribute ment_tsu8 of DEF_ARCH : architecture is " APB_PADDR[6]->APB_CLK=4.394";
   attribute ment_tsu9: string;
   attribute ment_tsu9 of DEF_ARCH : architecture is " APB_PADDR[7]->APB_CLK=4.459";
   attribute ment_tsu10: string;
   attribute ment_tsu10 of DEF_ARCH : architecture is " APB_PADDR[8]->APB_CLK=4.534";
   attribute ment_tsu11: string;
   attribute ment_tsu11 of DEF_ARCH : architecture is " APB_PADDR[9]->APB_CLK=4.111";
   attribute ment_tsu12: string;
   attribute ment_tsu12 of DEF_ARCH : architecture is " APB_PENABLE->APB_CLK=0.576";
   attribute ment_tsu13: string;
   attribute ment_tsu13 of DEF_ARCH : architecture is " APB_PSEL->APB_CLK=1.443";
   attribute ment_tsu14: string;
   attribute ment_tsu14 of DEF_ARCH : architecture is " APB_PWDATA[0]->APB_CLK=2.195";
   attribute ment_tsu15: string;
   attribute ment_tsu15 of DEF_ARCH : architecture is " APB_PWDATA[10]->APB_CLK=-0.156";
   attribute ment_tsu16: string;
   attribute ment_tsu16 of DEF_ARCH : architecture is " APB_PWDATA[11]->APB_CLK=-0.178";
   attribute ment_tsu17: string;
   attribute ment_tsu17 of DEF_ARCH : architecture is " APB_PWDATA[12]->APB_CLK=-0.110";
   attribute ment_tsu18: string;
   attribute ment_tsu18 of DEF_ARCH : architecture is " APB_PWDATA[13]->APB_CLK=-0.139";
   attribute ment_tsu19: string;
   attribute ment_tsu19 of DEF_ARCH : architecture is " APB_PWDATA[14]->APB_CLK=-0.131";
   attribute ment_tsu20: string;
   attribute ment_tsu20 of DEF_ARCH : architecture is " APB_PWDATA[15]->APB_CLK=-0.266";
   attribute ment_tsu21: string;
   attribute ment_tsu21 of DEF_ARCH : architecture is " APB_PWDATA[16]->APB_CLK=-0.048";
   attribute ment_tsu22: string;
   attribute ment_tsu22 of DEF_ARCH : architecture is " APB_PWDATA[17]->APB_CLK=-0.085";
   attribute ment_tsu23: string;
   attribute ment_tsu23 of DEF_ARCH : architecture is " APB_PWDATA[18]->APB_CLK=-0.079";
   attribute ment_tsu24: string;
   attribute ment_tsu24 of DEF_ARCH : architecture is " APB_PWDATA[19]->APB_CLK=-0.092";
   attribute ment_tsu25: string;
   attribute ment_tsu25 of DEF_ARCH : architecture is " APB_PWDATA[1]->APB_CLK=1.250";
   attribute ment_tsu26: string;
   attribute ment_tsu26 of DEF_ARCH : architecture is " APB_PWDATA[20]->APB_CLK=-0.052";
   attribute ment_tsu27: string;
   attribute ment_tsu27 of DEF_ARCH : architecture is " APB_PWDATA[21]->APB_CLK=-0.088";
   attribute ment_tsu28: string;
   attribute ment_tsu28 of DEF_ARCH : architecture is " APB_PWDATA[22]->APB_CLK=-0.108";
   attribute ment_tsu29: string;
   attribute ment_tsu29 of DEF_ARCH : architecture is " APB_PWDATA[23]->APB_CLK=-0.133";
   attribute ment_tsu30: string;
   attribute ment_tsu30 of DEF_ARCH : architecture is " APB_PWDATA[24]->APB_CLK=-0.076";
   attribute ment_tsu31: string;
   attribute ment_tsu31 of DEF_ARCH : architecture is " APB_PWDATA[25]->APB_CLK=-0.164";
   attribute ment_tsu32: string;
   attribute ment_tsu32 of DEF_ARCH : architecture is " APB_PWDATA[26]->APB_CLK=-0.256";
   attribute ment_tsu33: string;
   attribute ment_tsu33 of DEF_ARCH : architecture is " APB_PWDATA[27]->APB_CLK=-0.244";
   attribute ment_tsu34: string;
   attribute ment_tsu34 of DEF_ARCH : architecture is " APB_PWDATA[28]->APB_CLK=-0.134";
   attribute ment_tsu35: string;
   attribute ment_tsu35 of DEF_ARCH : architecture is " APB_PWDATA[29]->APB_CLK=-0.061";
   attribute ment_tsu36: string;
   attribute ment_tsu36 of DEF_ARCH : architecture is " APB_PWDATA[2]->APB_CLK=2.446";
   attribute ment_tsu37: string;
   attribute ment_tsu37 of DEF_ARCH : architecture is " APB_PWDATA[30]->APB_CLK=-0.080";
   attribute ment_tsu38: string;
   attribute ment_tsu38 of DEF_ARCH : architecture is " APB_PWDATA[31]->APB_CLK=-0.181";
   attribute ment_tsu39: string;
   attribute ment_tsu39 of DEF_ARCH : architecture is " APB_PWDATA[3]->APB_CLK=2.243";
   attribute ment_tsu40: string;
   attribute ment_tsu40 of DEF_ARCH : architecture is " APB_PWDATA[4]->APB_CLK=1.729";
   attribute ment_tsu41: string;
   attribute ment_tsu41 of DEF_ARCH : architecture is " APB_PWDATA[5]->APB_CLK=1.581";
   attribute ment_tsu42: string;
   attribute ment_tsu42 of DEF_ARCH : architecture is " APB_PWDATA[6]->APB_CLK=1.408";
   attribute ment_tsu43: string;
   attribute ment_tsu43 of DEF_ARCH : architecture is " APB_PWDATA[7]->APB_CLK=1.505";
   attribute ment_tsu44: string;
   attribute ment_tsu44 of DEF_ARCH : architecture is " APB_PWDATA[8]->APB_CLK=-0.161";
   attribute ment_tsu45: string;
   attribute ment_tsu45 of DEF_ARCH : architecture is " APB_PWDATA[9]->APB_CLK=-0.204";
   attribute ment_tsu46: string;
   attribute ment_tsu46 of DEF_ARCH : architecture is " APB_PWRITE->APB_CLK=1.482";
   attribute ment_tsu47: string;
   attribute ment_tsu47 of DEF_ARCH : architecture is " APB_RSTN->APB_CLK=2.569";
   attribute ment_tco0: string;
   attribute ment_tco0 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[0]=5.118";
   attribute ment_tco1: string;
   attribute ment_tco1 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[10]=4.443";
   attribute ment_tco2: string;
   attribute ment_tco2 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[11]=4.434";
   attribute ment_tco3: string;
   attribute ment_tco3 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[12]=4.433";
   attribute ment_tco4: string;
   attribute ment_tco4 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[13]=4.409";
   attribute ment_tco5: string;
   attribute ment_tco5 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[14]=4.407";
   attribute ment_tco6: string;
   attribute ment_tco6 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[15]=4.419";
   attribute ment_tco7: string;
   attribute ment_tco7 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[16]=4.423";
   attribute ment_tco8: string;
   attribute ment_tco8 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[17]=4.469";
   attribute ment_tco9: string;
   attribute ment_tco9 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[18]=4.438";
   attribute ment_tco10: string;
   attribute ment_tco10 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[19]=4.356";
   attribute ment_tco11: string;
   attribute ment_tco11 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[1]=5.053";
   attribute ment_tco12: string;
   attribute ment_tco12 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[20]=4.348";
   attribute ment_tco13: string;
   attribute ment_tco13 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[21]=4.716";
   attribute ment_tco14: string;
   attribute ment_tco14 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[22]=4.427";
   attribute ment_tco15: string;
   attribute ment_tco15 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[23]=4.654";
   attribute ment_tco16: string;
   attribute ment_tco16 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[24]=4.407";
   attribute ment_tco17: string;
   attribute ment_tco17 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[25]=4.369";
   attribute ment_tco18: string;
   attribute ment_tco18 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[26]=4.643";
   attribute ment_tco19: string;
   attribute ment_tco19 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[27]=4.484";
   attribute ment_tco20: string;
   attribute ment_tco20 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[28]=4.653";
   attribute ment_tco21: string;
   attribute ment_tco21 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[29]=4.235";
   attribute ment_tco22: string;
   attribute ment_tco22 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[2]=5.094";
   attribute ment_tco23: string;
   attribute ment_tco23 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[30]=4.499";
   attribute ment_tco24: string;
   attribute ment_tco24 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[31]=4.590";
   attribute ment_tco25: string;
   attribute ment_tco25 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[3]=4.851";
   attribute ment_tco26: string;
   attribute ment_tco26 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[4]=5.198";
   attribute ment_tco27: string;
   attribute ment_tco27 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[5]=5.068";
   attribute ment_tco28: string;
   attribute ment_tco28 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[6]=5.083";
   attribute ment_tco29: string;
   attribute ment_tco29 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[7]=5.613";
   attribute ment_tco30: string;
   attribute ment_tco30 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[8]=4.420";
   attribute ment_tco31: string;
   attribute ment_tco31 of DEF_ARCH : architecture is " APB_CLK->APB_PRDATA[9]=4.416";
   attribute ment_tco32: string;
   attribute ment_tco32 of DEF_ARCH : architecture is " APB_CLK->APB_PREADY=4.516";
   attribute ment_tco33: string;
   attribute ment_tco33 of DEF_ARCH : architecture is " APB_CLK->PCIE_SYSTEM_INT=3.967";
   attribute ment_tco34: string;
   attribute ment_tco34 of DEF_ARCH : architecture is " APB_CLK->PLL_LOCKLOST_INT=3.471";
   attribute ment_tco35: string;
   attribute ment_tco35 of DEF_ARCH : architecture is " APB_CLK->PLL_LOCK_INT=3.213";
   attribute ment_tco36: string;
   attribute ment_tco36 of DEF_ARCH : architecture is " REFCLK1->ATXCLKSTABLE[0]=2.210";
   attribute ment_tco37: string;
   attribute ment_tco37 of DEF_ARCH : architecture is " REFCLK1->ATXCLKSTABLE[1]=2.188";
   attribute black_box_pad : string;
   attribute black_box_pad of DEF_ARCH : architecture is "RXD3_P,RXD2_P,RXD1_P,RXD0_P,RXD3_N,RXD2_N,RXD1_N,RXD0_N,TXD3_P,TXD2_P,TXD1_P,TXD0_P,TXD3_N,TXD2_N,TXD1_N,TXD0_N";

begin

end DEF_ARCH;
