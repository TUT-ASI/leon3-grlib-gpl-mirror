-- Xilinx MIG Series 7
  constant CFG_MIG_SERIES7    : integer := CONFIG_MIG_SERIES7;
  constant CFG_MIG_SERIES7_MODEL    : integer := CONFIG_MIG_SERIES7_MODEL;

