
package version is
  constant grlib_version : integer := 2021100;
  constant grlib_build : integer := 4265;
end;
