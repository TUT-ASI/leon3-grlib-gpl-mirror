
package version is
  constant grlib_version : integer := 2023200;
  constant grlib_build : integer := 4283;
end;
