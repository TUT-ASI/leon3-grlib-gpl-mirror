-- High Speed Serial Links
  constant CFG_GRHSSL : integer := CONFIG_GRHSSL_ENABLE;
