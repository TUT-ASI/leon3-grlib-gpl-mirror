
package version is
  constant grlib_version : integer := 2018300;
  constant grlib_build : integer := 4226;
end;
