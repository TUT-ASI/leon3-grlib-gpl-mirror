
package version is
  constant grlib_version : integer := 2024100;
  constant grlib_build : integer := 4292;
end;
