
package version is
  constant grlib_version : integer := 2023400;
  constant grlib_build : integer := 4288;
end;
