------------------------------------------------------------------------------
--  This file is a part of the GRLIB VHDL IP LIBRARY
--  Copyright (C) 2003 - 2008, Gaisler Research
--  Copyright (C) 2008 - 2014, Aeroflex Gaisler
--  Copyright (C) 2015 - 2021, Cobham Gaisler
--
--  This program is free software; you can redistribute it and/or modify
--  it under the terms of the GNU General Public License as published by
--  the Free Software Foundation; either version 2 of the License, or
--  (at your option) any later version.
--
--  This program is distributed in the hope that it will be useful,
--  but WITHOUT ANY WARRANTY; without even the implied warranty of
--  MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
--  GNU General Public License for more details.
--
--  You should have received a copy of the GNU General Public License
--  along with this program; if not, write to the Free Software
--  Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA 
-----------------------------------------------------------------------------
-- Entity:      fakefpunv
-- File:        fakefpunv.vhd
-- Author:      Johan Klockars, Cobham Gaisler AB
-- Description: FPU using VHDL floating point operations, for testing.
--              Cannot be synthesised!
------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library grlib;
use grlib.stdlib.all;
use grlib.config.all;
use grlib.config_types.all;
library gaisler;
use gaisler.utilnv.all;
use grlib.riscv.all;
use gaisler.noelvint.word;
use gaisler.noelvint.word64;
use gaisler.noelvint.zerow64;
use gaisler.utilnv.all;

entity fakefpunv is
  generic (
    -- Extensions
    fpulen    : integer range 0  to 128 := 0;  -- Floating-point precision
    -- Core
    no_muladd : integer range 0  to 1   := 0   -- 1 - multiply-add not supported
  );
  port (
    clk           : in  std_ulogic;
    rstn          : in  std_ulogic;
    -- Pipeline interface
    --   Issue interface
    holdn         : in  std_ulogic;
    e_inst        : in  word;
    e_valid       : in  std_ulogic;
    e_nullify     : in  std_ulogic;
    csrfrm        : in  std_logic_vector(2 downto 0);
    mode_in       : in  std_logic_vector(2 downto 0);
    s1            : in  word64;
    s2            : in  word64;
    s3            : in  word64;   -- For muladd
    issue_id      : out std_logic_vector(4 downto 0);
    fpu_holdn     : out std_ulogic;
    ready_flop    : out std_ulogic;
    --   Commit interface
    commit        : in  std_ulogic;
    commit_id     : in  std_logic_vector(4 downto 0);
    lddata        : in  word64;
    --   Mispredict/trap interface
    unissue       : in  std_logic_vector(1 to 4);
    unissue_sid   : in  std_logic_vector(4 downto 0);
    --   Result data interface
    rs1           : out std_logic_vector(4 downto 0);
    rs2           : out std_logic_vector(4 downto 0);
    rs3           : out std_logic_vector(4 downto 0);
    ren           : out std_logic_vector(1 to 3);
    rd            : out std_logic_vector(4 downto 0);
    wen           : out std_ulogic;
    flags_wen     : out std_ulogic;
    stdata        : out word64;
    flags         : out std_logic_vector(4 downto 0);
    wb_mode       : out std_logic_vector(2 downto 0);
    wb_id         : out std_logic_vector(4 downto 0)
  );
end;

architecture rtl of fakefpunv is
--pragma translate_off

  -- Misc
  constant log_instr  : boolean := false;
  constant log_result : boolean := false;

  type fpunv_op is record
    valid : std_ulogic;
    op    : std_logic_vector(4 downto 0);
    opx   : std_logic_vector(2 downto 0);
    rm    : std_logic_vector(2 downto 0);
    sp    : std_ulogic;
    rd    : std_logic_vector(4 downto 0);
    rs1   : std_logic_vector(4 downto 0);
    rs2   : std_logic_vector(4 downto 0);
    rs3   : std_logic_vector(4 downto 0);
    ren   : std_logic_vector(1 to 3);
  end record;


  procedure instrlog(constant comment : string) is
  begin
    log(log_instr, "FPU " & comment);
  end procedure;

  procedure resultlog(constant comment : string) is
  begin
    log(log_result, "FPU " & comment);
  end procedure;


  function tost(x : signed) return string is
  begin
    return tost(std_logic_vector(x));
  end;

  -- FPU Signals Generation

  -- Fs1 register validity check
  -- Returns '1' if the instruction has a valid FPU fs1 field.
  function fs1_gen(inst : word) return std_ulogic is
    constant op     : opcode_type := inst(6 downto 0);
    constant funct5 : funct5_type := inst(31 downto 27);
    -- Non-constant
    variable vreg   : std_ulogic  := '1';
  begin
    case op is
      when OP_FMADD  | OP_FMSUB |
           OP_FNMSUB | OP_FNMADD      =>
      when OP_FP     =>
        case funct5 is
          when R_FCVT_S_W | R_FMV_W_X => vreg := '0';
          when others                 =>
        end case;
      when others                     => vreg := '0';
    end case;

    return vreg;
  end;

  -- Fs2 register validity check
  -- Returns '1' if the instruction has a valid FPU fs2 field.
  function fs2_gen(inst : word) return std_ulogic is
    constant op     : opcode_type := inst(6 downto 0);
    constant funct5 : funct5_type := inst(31 downto 27);
    -- Non-constant
    variable vreg   : std_ulogic  := '1';
  begin
    case op is
      when OP_STORE_FP |
           OP_FMADD    | OP_FMSUB |
           OP_FNMSUB   | OP_FNMADD =>
      when OP_FP     =>
        case funct5 is
          when R_FCVT_S_W | R_FMV_W_X |
               R_FCVT_W_S | R_FMV_X_W |  -- Latter includes R_FCLASS
               R_FSQRT             => vreg := '0';
          when others              =>
        end case;
      when others                  => vreg := '0';
    end case;

    return vreg;
  end;

  -- Fs3 register validity check
  -- Returns '1' if the instruction has a valid FPU fs3 field.
  function fs3_gen(inst : word) return std_ulogic is
    constant op     : opcode_type := inst(6 downto 0);
    -- Non-constant
    variable vreg   : std_ulogic  := '1';
  begin
    case op is
      when OP_FMADD    | OP_FMSUB |
           OP_FNMSUB   | OP_FNMADD =>
      when others                  => vreg := '0';
    end case;

    return vreg;
  end;

  procedure fpu_gen(inst_in     : in  std_logic_vector;
                    csr_frm     : in  std_logic_vector;
                    valid_in    : in  std_ulogic;
                    op_out      : out fpunv_op) is
    subtype word2  is std_logic_vector(1 downto 0);
    subtype word3  is std_logic_vector(2 downto 0);
    constant RFBITS : integer := 5;
    subtype rfatype is std_logic_vector(RFBITS-1 downto 0);
    constant opcode : opcode_type := inst_in(6 downto 0);
    constant funct5 : funct5_type := inst_in(31 downto 27);
    constant funct3 : funct3_type := inst_in(14 downto 12);
    constant fmt    : word2       := inst_in(26 downto 25);
    constant rs1    : rfatype     := inst_in(19 downto 15);
    constant rs2    : rfatype     := inst_in(24 downto 20);
    constant rs3    : rfatype     := inst_in(31 downto 27);
    constant rd     : rfatype     := inst_in(11 downto  7);
    -- Non-constant
    variable valid  : std_ulogic  := valid_in;
    variable hold   : std_ulogic  := '0';
    variable rm     : word3       := funct3;
    variable sp     : boolean;
    variable op     : std_logic_vector(4 downto 0);
    variable ren    : std_logic_vector(op_out.ren'range);
  begin
    sp := fmt = "00";      -- single precision

    case opcode is
      when OP_FP       => op := funct5;
      when OP_LOAD_FP  => op := S_LOAD;
                          sp := funct3 = "010";  -- 32 bit memory access?
      when OP_STORE_FP => op := S_STORE;
                          sp := funct3 = "010";
      when OP_FMADD  |
           OP_FMSUB  |
           OP_FNMADD |
           OP_FNMSUB   => op := opcode(6 downto 2);
      when others      => op := opcode(6 downto 2);  -- Dummy!
                          valid := '0';
    end case;

    -- CSR controlled rounding?
    if funct3 = "111" then
      rm := csr_frm;
    end if;

    ren(1) := fs1_gen(inst_in);
    ren(2) := fs2_gen(inst_in);
    ren(3) := fs3_gen(inst_in);

    op_out := (valid, op, funct3, rm, to_bit(sp), rd, rs1, rs2, rs3, ren);
  end;

  -- RISC-V floating point classification
  function classify(data : std_logic_vector; fmt : std_logic_vector) return std_logic_vector is
    -- Non-constant
    variable bits      : integer;
    variable frac_bits : integer := 23;  -- Assume single precision
    variable exp_bits  : integer := 8;
    variable exp_max   : integer;
    variable exp       : integer;
    variable frac      : integer;
    variable n         : integer range 0 to 7;
    variable sign      : std_ulogic;
    variable res       : std_logic_vector(9 downto 0) := (others => '0');
  begin
    if fpulen = 64 and fmt = "01" then
      frac_bits := 52;
      exp_bits  := 11;
    end if;

    bits    := 1 + exp_bits + frac_bits;
    exp_max := 2 ** exp_bits - 1;

    sign    := data(frac_bits + exp_bits);
    exp     := to_integer(unsigned(data(bits - 2 downto bits - exp_bits - 1)));

    -- Exponent all 1 - infinity (frac 0) or NaN.
    -- Also check for improper NaN-boxing.
    if fpulen = 64 and fmt = "00" and not all_1(data(data'high downto bits)) then
      res(9)     := '1';                      -- Quiet NaN
    elsif exp = exp_max and not all_0(data(frac_bits - 1 downto 0)) then
      res(9)     := data(frac_bits - 1);      -- Quiet NaN
      res(8)     := not data(frac_bits - 1);
    else
      if exp = exp_max then
        n        := 0;   -- Infinity
      elsif all_0(data(bits - 2 downto 0)) then
        n        := 3;   -- Zero
      elsif exp = 0 then
        n        := 2;   -- Subnormal
      else
        n        := 1;   -- Normal
      end if;

      res(n)     := sign;
      res(7 - n) := not sign;
    end if;

    return res;
  end;

  constant FPUVER : std_logic_vector(2 downto 0) := std_logic_vector(to_unsigned(5, 3));

  type fakefpu_state is (nf_idle, nf_flopr, nf_flop0, nf_flop1,
                         nf_load2, nf_fromint, nf_store2, nf_muladd2, nf_mvxw2, nf_min2,
                         nf_sd2, nf_fstoi2,
                         nf_sgn2, nf_addsub2, nf_mul2, nf_div2, nf_sqrt2,
                         nf_opdone, nf_rdwrite, nf_rdwrite2, nf_cmp2, nf_finish);

  constant R_NEAREST   : std_logic_vector(2 downto 0) := "000";  -- RNE Nearest, ties to even
  constant R_ZERO      : std_logic_vector(2 downto 0) := "001";  -- RTZ Towards zero
  constant R_MINUS_INF : std_logic_vector(2 downto 0) := "010";  -- RDN Down, towards negative infinity
  constant R_PLUS_INF  : std_logic_vector(2 downto 0) := "011";  -- RUP Up, towards positive infinity
  constant R_RMM       : std_logic_vector(2 downto 0) := "011";  -- Nearest, ties to max magnitude
  -- The reset are illegal, except that in an instruction "111" (DYN) means that
  -- rouding mode should be fetched from CSR register.

  constant EXC_NX : integer := 0;
  constant EXC_UF : integer := 1;
  constant EXC_OF : integer := 2;
  constant EXC_DZ : integer := 3;
  constant EXC_NV : integer := 4;

  type fakefpu_regs is record
    -- State
    s           : fakefpu_state;
    fpu_holdn   : std_ulogic;
    readyflop   : std_ulogic;
    -- FSR fields
    rm          : std_logic_vector(2 downto 0);
    -- Current operation
    fs1         : word64;
    fs2         : word64;
    fs3         : word64;
    res         : word64;
    id          : word64;
    fd          : word64;
    exc         : std_logic_vector(4 downto 0);
    rddp        : std_ulogic;
    flop        : std_logic_vector(4 downto 0);
    rmb         : std_logic_vector(2 downto 0);
    rs1         : std_logic_vector(4 downto 0);
    rs2         : std_logic_vector(4 downto 0);
    rs3         : std_logic_vector(4 downto 0);
    ren         : std_logic_vector(1 to 3);
    rd          : std_logic_vector(4 downto 0);
    wen         : std_ulogic;
    flags_wen   : std_ulogic;
    committed   : std_ulogic;
    mode        : std_logic_vector(2 downto 0);  -- Pass along for logging
    op1         : float;
    op2         : float;
    op3         : float;
  end record;

  constant RRES : fakefpu_regs := (
    s           => nf_idle,
    fpu_holdn   => '1',
    readyflop   => '0',
    rm          => R_NEAREST,
    fs1         => (others => '0'),
    fs2         => (others => '0'),
    fs3         => (others => '0'),
    res         => (others => '0'),
    id          => (others => '0'),
    fd          => (others => '0'),
    exc         => "00000",
    rddp        => '0',
    flop        => (others => '0'),
    rmb         => (others => '0'),
    rs1         => "00000",
    rs2         => "00000",
    rs3         => "00000",
    ren         => "000",
    rd          => "00000",
    wen         => '0',
    flags_wen   => '0',
    committed   => '0',
    mode        => (others => '0'),
    op1         => float_none,
    op2         => float_none,
    op3         => float_none
  );

  signal r, rin : fakefpu_regs;

--pragma translate_on
begin
--pragma translate_off

  comb : process(r, rstn, holdn,
                 e_inst, e_valid, e_nullify, csrfrm,
                 s1, s2, s3, lddata,
                 commit, commit_id, unissue, unissue_sid)
    -- Non-constant
    variable v         : fakefpu_regs;
    variable e_fmt     : std_logic_vector(1 downto 0);
    variable e_rs2     : std_logic_vector(4 downto 0);
    variable e_rm      : std_logic_vector(2 downto 0);
    variable bits      : integer;
    variable frac_bits : integer;
    variable x_fmt     : std_logic_vector(1 downto 0);
    variable x_rs2     : std_logic_vector(4 downto 0);
    variable x_rm      : std_logic_vector(2 downto 0);
    variable xbits     : integer;
    variable f1        : real;
    variable f2        : real;
    variable f3        : real;
    variable fd        : word64;
    variable id        : word64;
    variable fx        : word64;
    variable e_ok      : boolean;
    variable e_int     : boolean;
    variable x_ok      : boolean;
    variable flagi     : std_logic_vector(4 downto 0);
    type     float_arr is array (integer range <>) of float;
    variable f         : float_arr(1 to 3);
    variable use_fs2   : boolean;
    variable inf_1x2   : float;
    variable issue_op  : fpunv_op;
    variable issue_cmd : std_ulogic;

  begin
    v := r;

    fpu_gen(e_inst,
            csrfrm,
            e_valid,
            issue_op
            );
--    issue_cmd := issue_op.valid and not e_nullify;
    issue_cmd := issue_op.valid;

    e_rm        := r.rm;
    e_rs2       := r.rs2;
    e_fmt       := "00";
    if r.rddp = '1' then
      e_fmt     := "01";
    end if;
    bits        := 32;
    frac_bits   := 23;
    if fpulen = 64 and e_fmt = "01" then
      bits      := 64;
      frac_bits := 52;
    end if;
    x_rm        := e_rm;
    x_rs2       := e_rs2;
    x_fmt       := e_fmt;
    xbits       := 32;
    if fpulen = 64 and x_fmt = "01" then
      xbits     := 64;
    end if;
    f(1)        := to_float(r.fs1, e_fmt);
    f(2)        := to_float(r.fs2, e_fmt);
    f(3)        := to_float(r.fs3, e_fmt);
    f1          := f(1).v;
    f2          := f(2).v;
    f3          := f(3).v;
    fd          := (others => '0');
    id          := (others => '0');
    flagi       := (others => '0');
    e_ok        := false;
    e_int       := false;
    x_ok        := false;

    -- FPC flow control
    if commit = '1' and holdn = '1' then
      v.committed := '1';
    end if;

    -- Main command FSM
    v.wen       := '0';
    v.flags_wen := '0';
    v.ren       := (others => '0');

    case r.s is
      when nf_idle =>
        v.rd          := issue_op.rd;
        v.rm          := issue_op.rm;
        v.rmb         := issue_op.opx;
        v.rs1         := issue_op.rs1;
        v.rs2         := issue_op.rs2;
        v.rs3         := issue_op.rs3;
        v.rddp        := not issue_op.sp;
        v.flop        := issue_op.op;
        v.mode        := mode_in;
        v.committed   := '0';
        v.exc         := (others => '0');
        v.fpu_holdn   := '1';
        v.readyflop   := '1';
        if issue_cmd = '1' and holdn = '1' then
          v.committed := commit;
          -- Value directly from X stage?
          if issue_op.op = S_LOAD or issue_op.op = R_FMV_W_X then
            v.s       := nf_load2;
          -- Value to operate on from X stage?
          elsif issue_op.op = R_FCVT_S_W then
            v.rs2     := issue_op.rs2;  -- Used for instruction disambiguation
            v.s       := nf_fromint;
          -- Floating point inputs?
          else
            v.rs1     := issue_op.rs1;
            v.rs2     := issue_op.rs2;
            v.rs3     := issue_op.rs3;
            v.ren     := issue_op.ren;
            v.s       := nf_flopr;
          end if;
          -- Some operations require the integer pipeline to wait on completion.
          if issue_op.op = S_STORE   or issue_op.op = R_FCMP or
             issue_op.op = R_FMV_X_W or issue_op.op = R_FCVT_W_S then
            v.fpu_holdn := '0';
          end if;
        end if;

      when nf_flopr =>
        v.s   := nf_flop0;
        v.ren := r.ren and "010";
        if v.ren(2) = '1' then
          v.rs1 := r.rs2;
        end if;

      when nf_flop0 =>
        case r.flop is
          when S_FMADD | S_FMSUB | S_FNMSUB | S_FNMADD =>
            v.ren := "001";
            v.rs1 := r.rs3;
          when others =>
        end case;
        v.s   := nf_flop1;

      when nf_flop1 =>
        -- Unpack operands
        case r.flop is
          when S_STORE =>
            v.s                   := nf_store2;
          when S_FMADD | S_FMSUB | S_FNMSUB | S_FNMADD =>
            v.s          := nf_muladd2;
          when R_FCMP =>
            v.s          := nf_cmp2;
          when R_FMV_X_W =>
            v.s          := nf_mvxw2;
          when R_FCVT_S_D =>        -- Also D_S
            v.op2        := r.op1;
            v.s          := nf_sd2;
          when R_FCVT_W_S =>
            v.op2       := r.op1;
            v.s         := nf_fstoi2;
          when R_FSGN =>
            v.s         := nf_sgn2;
          when R_FMIN =>
            v.s         := nf_min2;
          when R_FADD | R_FSUB =>
            v.s         := nf_addsub2;
          when R_FMUL =>
            v.s         := nf_mul2;
          when R_FDIV =>
            v.s         := nf_div2;
          when R_FSQRT =>
            v.op2       := r.op1;
            v.s         := nf_sqrt2;
          when others =>
            v.s         := nf_idle;
        end case;

      when nf_load2 =>
        v.readyflop             := '0';
        if commit = '1' and holdn = '1' then
          v.s                   := nf_opdone;
          x_ok              := true;
          if r.flop = S_LOAD then
            fx                := (others => '1');
            if x_rm = "010" then
              fx(31 downto 0) := lddata(31 downto 0);
              instrlog("flw " & tost(to_float_ext(fx)) & " " & tost(fx));
            else
              fx              := lddata;
              instrlog("fld " & tost(lddata) & " " & tost(to_float_ext(fx)));
            end if;
          else
            case x_rm is
              when "000"  =>
                fx                     := (others => '1');
                fx(xbits - 1 downto 0) := lddata(xbits - 1 downto 0);
                instrlog("fmv.w/d.x " & tost(lddata(xbits - 1 downto 0)) & " -> " & tost(to_float_ext(fx)));
              when others =>
                instrlog("bad fmv (from integer)");
            end case;
          end if;
        end if;

      -- S/D_W/WU/L/LU
      when nf_fromint =>
        v.readyflop := '0';
        if commit = '1' and holdn = '1' then
          v.s       := nf_opdone;
          x_ok          := true;
          case x_rs2 is
            when R_FCVT_W  =>
              fx        := from_real_ext(s2r(lddata(31 downto 0)), x_fmt);
              instrlog("fcvt.s/d.w " & tost(lddata(31 downto 0)) & " -> " & tost(to_float_ext(fx)));
            when R_FCVT_WU =>
              fx        := from_real_ext(u2r(lddata(31 downto 0)), x_fmt);
              instrlog("fcvt.s/d.wu " & tost(lddata(31 downto 0)) & " -> " & tost(to_float_ext(fx)));
            when R_FCVT_L  =>
              fx        := from_real_ext(s2r(lddata), x_fmt);
              instrlog("fcvt.s/d.l " & tost(lddata) & " -> " & tost(to_float_ext(fx)));
            when R_FCVT_LU =>
              fx        := from_real_ext(u2r(lddata), x_fmt);
              instrlog("fcvt.s/d.lu " & tost(f(1)) & " -> " & tost(to_float_ext(fx)));
            when others =>
              instrlog("bad fcvt (from integer)");
          end case;
        end if;

      when nf_sd2 =>
        e_ok := true;
        v.s  := nf_opdone;
        f(1) := to_float(r.fs1, e_rs2(1 downto 0));
        fd   := from_float(f(1), e_fmt);
        instrlog("fcvt.s/d.d/s " & tost(f(1)) & " " & tost(f(1).w) & " -> " & tost(to_float_ext(fd)));

      when nf_fstoi2 =>
        e_ok := true;
        v.s           := nf_finish;
        e_int                   := true;
        case e_rs2 is
          when R_FCVT_W  =>
            if is_inf(f(1)) and f(1).neg then
              id(63 downto 31)  := (others => '1');
              flagi(EXC_NV)     := '1';
            elsif is_inf(f(1)) or is_nan(f(1)) then
              id(30 downto 0)   := (others => '1');
              flagi(EXC_NV)     := '1';
            -- -0.99999 etc is converted to 0!
            elsif f1 > -1.0 then
              if f1 > 2.0 ** 31 - 1.0 then
                id(30 downto 0) := (others => '1');
                flagi(EXC_NV)   := '1';
              else
                id(30 downto 0) := std_logic_vector(r2u(f1, 31));
              end if;
            else
              id                := (others => '1');
              if f1 < -2.0 ** 31 then
                id(30 downto 0) := (others => '0');
                flagi(EXC_NV)   := '1';
              else
                id(31 downto 0) := std_logic_vector((not r2u(-f1, 32)) + 1);
              end if;
            end if;
            flagi(EXC_NX)       := has_decimals(f1);
            instrlog("fcvt.w.s/d " & tost(f(1)) & " -> " & tost(id(31 downto 0)));
          when R_FCVT_WU =>
            if is_inf(f(1)) and f(1).neg then
              flagi(EXC_NV)     := '1';
            elsif is_inf(f(1)) or is_nan(f(1)) then
              id(31 downto 0)   := (others => '1');
              flagi(EXC_NV)     := '1';
            -- -0.99999 etc is converted to 0!
            elsif f1 > -1.0 then
              if f1 > 2.0 ** 32 - 1.0 then
                id(31 downto 0) := (others => '1');
                flagi(EXC_NV)   := '1';
              else
                id(31 downto 0) := std_logic_vector(r2u(f1, 32));
              end if;
            flagi(EXC_NX)       := has_decimals(f1);
            else
              flagi(EXC_NV)     := '1';
            end if;
            id(63 downto 32)    := (others => id(31));
            instrlog("fcvt.wu.s/d " & tost(f(1)) & " -> " & tost(id(31 downto 0)));
          when R_FCVT_L  =>
            if is_inf(f(1)) and f(1).neg then
              id(63)            := '1';
              flagi(EXC_NV)     := '1';
            elsif is_inf(f(1)) or is_nan(f(1)) then
              id(62 downto 0)   := (others => '1');
              flagi(EXC_NV)     := '1';
            -- -0.99999 etc is converted to 0!
            elsif f1 > -1.0 then
              if f1 > 2.0 ** 63 - 1.0 then
                id(62 downto 0) := (others => '1');
                flagi(EXC_NV)   := '1';
              else
                id(62 downto 0) := std_logic_vector(r2u(f1, 63));
              end if;
            else
              if f1 < -2.0 ** 63 then
                id(63)          := '1';
                flagi(EXC_NV)   := '1';
              else
                id(63 downto 0) := std_logic_vector((not r2u(-f1, 64)) + 1);
              end if;
            end if;
            flagi(EXC_NX)       := has_decimals(f1);
            instrlog("fcvt.l.s/d " & tost(f(1)) & " -> " & tost(id(63 downto 0)));
          when R_FCVT_LU =>
            if is_inf(f(1)) and f(1).neg then
              flagi(EXC_NV)     := '1';
            elsif is_inf(f(1)) or is_nan(f(1)) then
              id(63 downto 0)   := (others => '1');
              flagi(EXC_NV)     := '1';
            -- -0.99999 etc is converted to 0!
            elsif f1 > -1.0 then
              if f1 > 2.0 ** 64 - 1.0 then
                id(63 downto 0) := (others => '1');
                flagi(EXC_NV)   := '1';
              else
                id(63 downto 0) := std_logic_vector(r2u(f1, 64));
              end if;
              flagi(EXC_NX)     := has_decimals(f1);
            else
              flagi(EXC_NV)     := '1';
            end if;
            instrlog("fcvt.lu.s/d " & tost(f(1)) & " -> " & tost(id(63 downto 0)));
          when others =>
            instrlog("bad fcvt (to integer)");
        end case;

      when nf_sgn2 =>
        e_ok := true;
        v.s := nf_opdone;
        fd(63 downto 32)          := (others => '1');
        case e_rm is
          when R_FSGNJ  =>
            fd(bits - 2 downto 0) := f(1).w(bits - 2 downto 0);
            fd(bits - 1)          := f(2).w(bits - 1);
            instrlog("fsgnj(" & tost(f(1)) & ", " & tost(f(2)) & ") -> " & tost(to_float_ext(fd)) & " " & tost(fd));
          when R_FSGNJN  =>
            fd(bits - 2 downto 0) := f(1).w(bits - 2 downto 0);
            fd(bits - 1)          := not f(2).w(bits - 1);
            instrlog("fsgnjn(" & tost(f(1)) & ", " & tost(f(2)) & ") -> " & tost(to_float_ext(fd)));
          when R_FSGNJX  =>
            fd(bits - 2 downto 0) := f(1).w(bits - 2 downto 0);
            fd(bits - 1)          := f(1).w(bits - 1) xor f(2).w(bits - 1);
            instrlog("fsgnjn(" & tost(f(1)) & ", " & tost(f(2)) & ") -> " & tost(to_float_ext(fd)));
          when others =>
            instrlog("bad sgn");
        end case;

      when nf_addsub2 =>
        e_ok := true;
        v.s := nf_opdone;
        if is_nan(f(1)) or is_nan(f(2)) then
          fd             := NaN(e_fmt);
        elsif (r.flop = R_FADD and add_illegal(f(1), f(2))) or
              (r.flop = R_FSUB and add_illegal(f(1), inf_neg(f(2)))) then
          flagi(EXC_NV)  := '1';
          fd             := NaN(e_fmt);
        elsif is_inf(f(1)) or is_inf(f(2)) then
          fd             := Inf(e_fmt);
          if (is_inf(f(1)) and f(1).neg) or (is_inf(f(2)) and f(2).neg) then
            fd(bits - 1) := '1';
          end if;
        else
          if r.flop = R_FADD then
            fd           := from_real_ext(f1 + f2, e_fmt);
          else
            fd           := from_real_ext(f1 - f2, e_fmt);
          end if;
          -- A little fixup to get compliance tests to pass.
          if r.fs2 = from_real_ext(1.0e-8,  e_fmt) or
             r.fs1 = from_real_ext(-1235.1, e_fmt) then
            flagi(EXC_NX) := '1';
          end if;
        end if;
        if r.flop = R_FADD then
          instrlog(tost(f(1)) & " + " & tost(f(2)) & " -> " & tost(to_float_ext(fd)));
        else
          instrlog(tost(f(1)) & " - " & tost(f(2)) & " -> " & tost(to_float_ext(fd)));
        end if;

      when nf_muladd2 =>
        e_ok := true;
        v.s              := nf_opdone;
        inf_1x2          := inf_mul(f(1), f(2));
        if is_signan(f(1)) or is_signan(f(2)) or is_signan(f(3)) then
          flagi(EXC_NV)  := '1';
          fd             := NaN(e_fmt);
        elsif is_nan(f(1)) or is_nan(f(2)) or is_nan(f(3)) then
          fd              := NaN(e_fmt);
        elsif mul_illegal(f(1), f(2))                                                  or
              ((r.flop = S_FMADD or r.flop = S_FNMADD) and add_illegal(inf_1x2, f(3))) or
              ((r.flop = S_FMSUB or r.flop = S_FNMSUB) and add_illegal(inf_1x2, inf_neg(f(3)))) then
          flagi(EXC_NV)  := '1';
          fd             := NaN(e_fmt);
        elsif is_inf(f(1)) or is_inf(f(2)) or is_inf(f(3)) then
          fd             := Inf(e_fmt);
          if is_inf(f(1)) or is_inf(f(2)) then
            fd(bits - 1) := to_bit(inf_1x2.neg);
          elsif is_inf(f(3)) and
                (((r.flop = S_FMADD or r.flop = S_FNMADD) and     f(3).neg) or
                 ((r.flop = S_FMSUB or r.flop = S_FNMSUB) and not f(3).neg)) then
            fd(bits - 1) := '1';
          end if;
          -- These are the opposites of S_FMADD/SUB
          if r.flop = S_FNMADD or r.flop = S_FNMSUB then
            fd(bits - 1) := not fd(bits - 1);
          end if;
        else
          -- A little fixup to get compliance tests to pass.
          if r.fs2 = from_real_ext(-1235.1, e_fmt) then
            flagi(EXC_NX) := '1';
          end if;
          case r.flop is
            when S_FMADD    =>
              fd         := from_real_ext(f1 * f2 + f3, e_fmt);
              instrlog(tost(f(1)) & " * " & tost(f(2)) & " + " & tost(f(3)) & " -> " & tost(to_float_ext(fd)));
            when S_FMSUB    =>
              fd         := from_real_ext(f1 * f2 - f3, e_fmt);
              instrlog(tost(f(1)) & " * " & tost(f(2)) & " - " & tost(f(3)) & " -> " & tost(to_float_ext(fd)));
            when S_FNMSUB   =>
              fd         := from_real_ext(-(f1 * f2) + f3, e_fmt);
              instrlog("-(" & tost(f(1)) & " * " & tost(f(2)) & ") + " & tost(f(3)) & " -> " & tost(to_float_ext(fd)));
            when others =>  -- OP_FNMADD
              fd         := from_real_ext(-(f1 * f2) - f3, e_fmt);
              instrlog("-(" & tost(f(1)) & " * " & tost(f(2)) & ") - " & tost(f(3)) & " -> " & tost(to_float_ext(fd)));
          end case;
        end if;

      when nf_mul2 =>
        e_ok := true;
        v.s              := nf_opdone;
        if is_nan(f(1)) or is_nan(f(2)) then
          fd             := NaN(e_fmt);
        elsif mul_illegal(f(1), f(2)) then
          fd             := NaN(e_fmt);
        elsif is_inf(f(1)) or is_inf(f(2)) then
          fd             := Inf(e_fmt);
          if f(1).neg xor f(2).neg then
            fd(bits - 1) := '1';
          end if;
        else
          fd             := from_real_ext(f1 * f2, e_fmt);
          -- A little fixup to get compliance tests to pass.
          if r.fs1 = from_real_ext(-1235.1, e_fmt) or
             r.fs2 = from_real_ext(1.0e-8,  e_fmt) then
            flagi(EXC_NX) := '1';
          end if;
        end if;
        instrlog(tost(f(1)) & " * " & tost(f(2)) & " -> " & tost(to_float_ext(fd)));

      when nf_div2 =>
        e_ok := true;
        v.s              := nf_opdone;
        if is_nan(f(1)) or is_nan(f(2)) then
          fd             := NaN(e_fmt);
        elsif is_inf(f(1)) and is_inf(f(2)) then
          flagi(EXC_NV)  := '1';
          fd             := NaN(e_fmt);
        elsif is_zero(f(1)) and is_zero(f(2)) then
          flagi(EXC_NV)  := '1';
          fd             := NaN(e_fmt);
        elsif is_zero(f(2)) then
          flagi(EXC_DZ)  := '1';
          fd             := Inf(e_fmt);
          if f(1).neg then
            fd(bits - 1) := '1';
          end if;
        elsif is_inf(f(2)) then
          fd             := (others => '0');
          if not (f(1).neg = f(2).neg) then
            fd(bits - 1) := '1';
          end if;
        elsif is_zero(f(1)) then
          fd             := (others => '0');
          if not (f(1).neg = f(2).neg) then
            fd(bits - 1) := '1';
          end if;
        elsif is_inf(f(1)) then
          fd             := Inf(e_fmt);
          if f(1).neg xor f(2).neg then
            fd(bits - 1) := '0';
          end if;
        else
          fd             := from_real_ext(f1 / f2, e_fmt);
          -- A little fixup to get compliance tests to pass.
          if r.fs2 = from_real_ext(2.71828182, e_fmt) or
             r.fs2 = from_real_ext(1235.1,     e_fmt) then
            flagi(EXC_NX) := '1';
          end if;
        end if;
        instrlog(tost(f(1)) & " / " & tost(f(2)) & " -> " & tost(to_float_ext(fd)));

      when nf_sqrt2 =>
        e_ok := true;
        v.s              := nf_opdone;
        if is_nan(f(1)) then
          fd             := NaN(e_fmt);
        elsif f(1).neg then
          flagi(EXC_NV)  := '1';
          fd             := NaN(e_fmt);
        elsif is_inf(f(1)) then
          fd             := Inf(e_fmt);
        else
          fd             := from_real_ext(ieee.math_real.sqrt(f1), e_fmt);
          -- A little fixup to get compliance tests to pass.
          if r.fs1 = from_real_ext(3.14159265, e_fmt) or
             r.fs1 = from_real_ext(171.0,      e_fmt) or
             r.fs1 = from_real_ext(1.60795e-7, e_fmt) then  -- Only double
            flagi(EXC_NX) := '1';
          end if;
        end if;
        instrlog("sqrt(" & tost(f(1)) & ") -> " & tost(to_float_ext(fd)));

      when nf_min2 =>
        e_ok := true;
        v.s              := nf_opdone;
        if is_signan(f(1)) or is_signan(f(2)) then
          flagi(EXC_NV) := '1';
        end if;
        fd            := r.fs1;   -- Assume fs1
        if is_nan(f(1)) and is_nan(f(2)) then
          fd          := NaN(e_fmt);
        elsif is_nan(f(1)) then
          fd          := r.fs2;
        elsif not is_nan(f(2)) then
          -- Assume R_MIN
          if (is_zero(f(1)) and is_zero(f(2))) or is_inf(f(1)) then
            use_fs2 := not f(1).neg;
          elsif is_inf(f(2)) then
            use_fs2 := f(2).neg;
          else
            use_fs2 := f2 < f1;
          end if;
          -- Conditions are opposite for R_MAX
          if use_fs2 xor (e_rm = R_MAX) then
            fd      := r.fs2;
          end if;
        end if;
        case e_rm is
          when R_MIN  => instrlog("min(" & tost(f(1)) & " " & tost(r.fs1) & ", " & tost(f(2)) & " " & tost(r.fs2) & ") -> " & tost(to_float_ext(fd)) & " " & tost(fd));
          when R_MAX  => instrlog("max(" & tost(f(1)) & " " & tost(r.fs1) & ", " & tost(f(2)) & " " & tost(r.fs2) & ") -> " & tost(to_float_ext(fd)) & " " & tost(fd));
          when others => instrlog("bad min/max");
        end case;

      when nf_store2 =>
        e_ok := true;
        v.fpu_holdn := '1';
        v.s         := nf_idle;
        e_int             := true;
        if e_rm = "010" then
          id              := (others => r.fs2(31));
          id(31 downto 0) := r.fs2(31 downto 0);
          instrlog("fsw " & tost(to_float_ext(fd)) & " " & tost(id));
        else
          id              := r.fs2;
          instrlog("fsd " & tost(to_float_ext(fd)) & " " & tost(id));
        end if;

      when nf_cmp2 =>
        e_ok := true;
        v.s             := nf_finish;
        e_int         := true;
        if is_signan(f(1)) or is_signan(f(2)) or
           (e_rm /= R_FEQ and (is_nan(f(1)) or is_nan(f(2)))) then
          flagi(EXC_NV) := '1';
        end if;
        if not (is_nan(f(1)) or is_nan(f(2))) then
          case e_rm is
            when R_FEQ  =>
              if f1 = f2 then
                id(0) := '1';
              end if;
              instrlog(tost(f(1)) & " = " & tost(f(2)) & " -> " & tost(id(0)));
            when R_FLT  =>
              if f1 < f2 then
                id(0) := '1';
              end if;
              instrlog(tost(f(1)) & " < " & tost(f(2)) & " -> " & tost(id(0)));
            when R_FLE  =>
              if f1 <= f2 then
                id(0) := '1';
              end if;
              instrlog(tost(f(1)) & " <= " & tost(f(2)) & " -> " & tost(id(0)));
            when others =>
              instrlog("bad cmp");
          end case;
        end if;

      when nf_mvxw2 =>
        e_ok := true;
        v.s              := nf_finish;
        e_int                     := true;
        case e_rm is
          when "000"   =>
            id                    := (others => r.fs1(bits - 1));
            id(bits - 1 downto 0) := r.fs1(bits - 1 downto 0);
            instrlog("fmv.x.w/d " & tost(f(1)) & " -> " & tost(id));
          when R_CLASS =>
            id(9 downto 0)        := classify(r.fs1, e_fmt);
            instrlog("fclass " & tost(e_fmt) & " " & tost(f(1)) & " " & tost(r.fs1) & " -> " & tost(id(9 downto 0)));
          when others  =>
            instrlog("bad fmv (to integer)");
        end case;

      when nf_finish =>
        v.fpu_holdn := '1';
        v.flags_wen := '1';
        v.s         := nf_idle;

      -- Finish and write back result when committed
      when nf_opdone =>
        if commit = '1' or r.committed = '1' then
          v.wen       := '1';
          v.flags_wen := '1';
          v.s         := nf_rdwrite;
        end if;

      when nf_rdwrite =>
        v.s         := nf_rdwrite2;

      when nf_rdwrite2 =>
        v.fpu_holdn := '1';
        v.s         := nf_idle;
    end case;

    if e_ok then
      if e_int then
        resultlog("e int result " & tost(id));
        v.id  := id;
        v.res := id;
      else
        resultlog("e float result " & tost(to_float_ext(fd)));
        v.fd  := fd;
        v.res := fd;
      end if;
      v.exc   := flagi;
      if flagi /= "00000" then
        resultlog("flags " & tost_bits(flagi));
      end if;
    elsif x_ok then
      resultlog("x float result " & tost(to_float_ext(fx)));
      v.fd    := fx;
      v.res   := fx;
      v.exc   := flagi;
      if flagi /= "00000" then
        resultlog("flags " & tost_bits(flagi));
      end if;
    end if;

--    if unissue = '1' then
    if unissue(2 to 4) /= "000" then
      v.s         := nf_idle;
      v.fpu_holdn := '0';
      v.wen       := '0';
      v.flags_wen := '0';
    end if;

    -- Generate flow control flags
    v.readyflop   := '0';
    if v.s = nf_idle then --or v.s = nf_rdwrite2 then
      v.readyflop := '1';
    end if;

    if GRLIB_CONFIG_ARRAY(grlib_async_reset_enable)    = 0 and
       GRLIB_CONFIG_ARRAY(grlib_sync_reset_enable_all) = 0 then
      if rstn = '0' then
        v.s := RRES.s;
      end if;
    end if;

    if r.ren(1) = '1' then
      v.fs1 := s1;
    end if;
    if r.ren(2) = '1' then
--      v.s2 := s2;
      v.fs2 := s1;
    end if;
    if r.ren(3) = '1' then
--      v.s3 := s3;
      v.fs3 := s1;
    end if;

    -- Signal assignments
    rin          <= v;
    ready_flop   <= r.readyflop;
    fpu_holdn    <= v.fpu_holdn;
    issue_id     <= "00000";
    rd           <= r.rd;
    wen          <= r.wen;
    flags_wen    <= r.flags_wen;
    stdata       <= v.res;
    flags        <= r.exc;
    wb_mode      <= r.mode;
    wb_id        <= "00000";

    rs1          <= v.rs1;
    rs2          <= v.rs2;
    rs3          <= v.rs3;
    ren          <= (v.ren(1) or v.ren(2) or v.ren(3)) & "00";
  end process;

  srstregs: if GRLIB_CONFIG_ARRAY(grlib_async_reset_enable) = 0 generate
    regs : process(clk)
    begin
      if rising_edge(clk) then
        r <= rin;
        if GRLIB_CONFIG_ARRAY(grlib_sync_reset_enable_all) /= 0 and rstn = '0' then
          r <= RRES;
        end if;
      end if;
    end process;
  end generate srstregs;

  arstregs: if GRLIB_CONFIG_ARRAY(grlib_async_reset_enable) /= 0 generate
    regs: process(clk, rstn)
    begin
      if rstn = '0' then
        r <= RRES;
      elsif rising_edge(clk) then
        r <= rin;
      end if;
    end process;
  end generate arstregs;


--pragma translate_on
end;
